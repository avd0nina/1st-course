`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 21.03.2024 03:13:49
// Design Name: 
// Module Name: count4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module count4(
    input clk,
    input lever,
    output logic [3:0] q
    );
    always_ff @(posedge clk) begin
//      q[0] <= !q[0];
//      q[1] <= q[1] ^ q[0];
//      q[2] <= q[2] ^ (q[1] & q[0]);
//      q <= q + 1;

//        q[0] <= !q[2] & !q[1] & !q[0]
//            | !q[2] & q[1] & !q[0];
//        q[1] <= !q[2] & !q[1] & q[0]
//            | !q[2] & q[1] & !q[0];
//        q[2] <= !q[2] & q[1] & q[0];

//        q[0] <= !q[0];
//        q[1] <= q[1] ^ ((!q[0] & !lever)
//                | (q[0] & lever));
//        q[2] <= q[2] ^ (((!q[1] & !q[0]) & !lever)
//        | ((q[1] & q[0]) & lever));
//        q[3] <= q[3] ^ (((!q[2] & !q[1] & !q[0]) & !lever)
//        | ((q[2] & q[1] & q[0]) & lever));

//        q[0] <= !q[0] & !q[1] & !q[2] & !q[3]
//            | !q[0] & q[1] & !q[2] & !q[3]
//            | !q[0] & !q[1] & q[2] & !q[3]
//            | !q[0] & q[1] & q[2] & !q[3]
//            | !q[0] & !q[1] & !q[2] & q[3]
//            | !q[0] & q[1] & !q[2] & q[3];
            
        q[0] <= !q[0];
        
        q[1] <= (lever & (q[0] & !q[1] & !q[2] & !q[3]
            | !q[0] & q[1] & !q[2] & !q[3]
            | q[0] & !q[1] & q[2] & !q[3]
            | !q[0] & q[1] & q[2] & !q[3]
            | q[0] & !q[1] & !q[2] & q[3]
            | !q[0] & q[1] & !q[2] & q[3]))
        | (!lever & (!q[0] & !q[1] & !q[2] & !q[3]
            | q[0] & q[1] & !q[2] & !q[3]
            | !q[0] & !q[1] & q[2] & !q[3]
            | q[0] & q[1] & q[2] & !q[3]
            | !q[0] & !q[1] & !q[2] & q[3]
            | q[0] & q[1] & !q[2] & q[3]));
        
        q[2] <= (lever & (q[0] & q[1] & !q[2] & !q[3]
            | !q[0] & !q[1] & q[2] & !q[3]
            | q[0] & !q[1] & q[2] & !q[3]
            | !q[0] & q[1] & q[2] & !q[3]))
        | (!lever & (q[0] & !q[1] & q[2] & !q[3]
            | !q[0] & q[1] & q[2] & !q[3]
            | q[0] & q[1] & q[2] & !q[3]
            | !q[0] & !q[1] & !q[2] & q[3]));
        
        q[3] <= (lever & (q[0] & q[1] & q[2] & !q[3]
            | !q[0] & !q[1] & !q[2] & q[3]
            | q[0] & !q[1] & !q[2] & q[3]
            | !q[0] & q[1] & !q[2] & q[3]))
         | (!lever & (!q[0] & !q[1] & !q[2] & !q[3]
            | q[0] & !q[1] & !q[2] & q[3]
            | !q[0] & q[1] & !q[2] & q[3]
            | q[0] & q[1] & !q[2] & q[3]));
   end
endmodule
